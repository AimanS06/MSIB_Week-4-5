magic
tech sky130A
magscale 1 2
timestamp 1729412534
<< nwell >>
rect -217 -1748 655 679
<< nsubdiff >>
rect -181 609 -121 643
rect 559 609 619 643
rect -181 583 -147 609
rect 585 583 619 609
rect -181 -1678 -147 -1652
rect 585 -1678 619 -1652
rect -181 -1712 -121 -1678
rect 559 -1712 619 -1678
<< nsubdiffcont >>
rect -121 609 559 643
rect -181 -1652 -147 583
rect 585 -1652 619 583
rect -121 -1712 559 -1678
<< poly >>
rect 6 69 36 111
rect -57 53 36 69
rect -57 19 -41 53
rect -7 19 36 53
rect -57 3 36 19
rect 6 2 36 3
rect 410 69 440 79
rect 410 53 502 69
rect 410 19 452 53
rect 486 19 502 53
rect 410 3 502 19
rect 410 2 440 3
rect 5 -444 36 -409
rect -56 -460 36 -444
rect -56 -494 -40 -460
rect -6 -494 36 -460
rect 410 -435 440 -393
rect 410 -451 501 -435
rect -56 -510 36 -494
rect 93 -594 193 -480
rect 252 -591 351 -483
rect 410 -485 451 -451
rect 485 -485 501 -451
rect 410 -501 501 -485
rect 410 -502 440 -501
rect 409 -565 501 -549
rect 409 -599 451 -565
rect 485 -599 501 -565
rect 409 -615 501 -599
rect 409 -660 439 -615
rect 5 -927 35 -901
rect -58 -943 35 -927
rect -58 -977 -42 -943
rect -8 -977 35 -943
rect -58 -993 35 -977
rect -58 -1096 35 -1080
rect -58 -1130 -42 -1096
rect -8 -1130 35 -1096
rect -58 -1146 35 -1130
rect 4 -1153 35 -1146
rect 408 -1096 500 -1080
rect 408 -1130 450 -1096
rect 484 -1130 500 -1096
rect 408 -1146 500 -1130
rect 408 -1154 438 -1146
<< polycont >>
rect -41 19 -7 53
rect 452 19 486 53
rect -40 -494 -6 -460
rect 451 -485 485 -451
rect 451 -599 485 -565
rect -42 -977 -8 -943
rect -42 -1130 -8 -1096
rect 450 -1130 484 -1096
<< locali >>
rect -181 609 -121 643
rect 559 609 619 643
rect -181 583 -147 609
rect 585 583 619 609
rect -57 19 -41 53
rect -7 19 9 53
rect 436 19 452 53
rect 486 19 502 53
rect -56 -494 -40 -460
rect -6 -494 10 -460
rect 435 -485 451 -451
rect 485 -485 501 -451
rect 435 -599 451 -565
rect 485 -599 501 -565
rect -58 -977 -42 -943
rect -8 -977 8 -943
rect -58 -1130 -42 -1096
rect -8 -1130 8 -1096
rect 434 -1130 450 -1096
rect 484 -1130 500 -1096
rect -181 -1678 -147 -1652
rect 585 -1678 619 -1652
rect -181 -1712 -121 -1678
rect 559 -1712 619 -1678
<< viali >>
rect 68 609 199 643
rect -41 19 -7 53
rect 452 19 486 53
rect -40 -494 -6 -460
rect 451 -485 485 -451
rect 451 -599 485 -565
rect -42 -977 -8 -943
rect -42 -1130 -8 -1096
rect 450 -1130 484 -1096
<< metal1 >>
rect 56 643 211 649
rect 56 609 68 643
rect 199 609 211 643
rect 56 603 211 609
rect 444 554 454 560
rect 0 513 454 554
rect 0 300 43 513
rect 444 508 454 513
rect 506 508 516 560
rect -52 100 94 300
rect 187 176 197 228
rect 249 176 259 228
rect 352 100 399 300
rect 451 100 498 300
rect -41 59 -6 100
rect -53 53 5 59
rect -53 19 -41 53
rect -7 19 5 53
rect -53 13 5 19
rect 123 -22 165 53
rect 266 10 276 62
rect 328 10 338 62
rect 452 59 486 100
rect 440 53 498 59
rect 440 19 452 53
rect 486 19 498 53
rect 440 13 498 19
rect 123 -64 322 -22
rect 106 -154 116 -102
rect 168 -154 178 -102
rect 280 -146 322 -64
rect -59 -393 -49 -193
rect 3 -393 94 -193
rect 352 -267 498 -193
rect 185 -322 195 -267
rect 252 -322 262 -267
rect 352 -323 441 -267
rect 497 -323 507 -267
rect 352 -393 498 -323
rect -40 -454 -6 -393
rect 439 -451 497 -393
rect -52 -460 6 -454
rect -52 -494 -40 -460
rect -6 -494 6 -460
rect 439 -485 451 -451
rect 485 -485 497 -451
rect 439 -491 497 -485
rect -52 -500 6 -494
rect 439 -565 497 -559
rect 439 -599 451 -565
rect 485 -599 497 -565
rect -60 -885 -50 -685
rect 2 -885 93 -685
rect 439 -686 497 -599
rect 351 -762 497 -686
rect 183 -822 193 -764
rect 251 -822 261 -764
rect 351 -818 440 -762
rect 496 -818 506 -762
rect -42 -937 -6 -885
rect 351 -886 497 -818
rect -54 -943 4 -937
rect -54 -977 -42 -943
rect -8 -977 4 -943
rect 106 -975 116 -923
rect 168 -975 178 -923
rect -54 -983 4 -977
rect 282 -1004 321 -932
rect 123 -1043 321 -1004
rect -54 -1096 4 -1090
rect -54 -1130 -42 -1096
rect -8 -1130 4 -1096
rect 123 -1130 162 -1043
rect -54 -1136 4 -1130
rect -42 -1177 -7 -1136
rect 264 -1139 274 -1087
rect 326 -1139 336 -1087
rect 438 -1096 496 -1090
rect 438 -1130 450 -1096
rect 484 -1130 496 -1096
rect 438 -1136 496 -1130
rect 450 -1177 484 -1136
rect -54 -1377 92 -1177
rect 183 -1305 193 -1247
rect 251 -1305 261 -1247
rect 350 -1377 397 -1177
rect 449 -1377 496 -1177
rect -2 -1568 40 -1377
rect 445 -1562 455 -1556
rect 442 -1568 455 -1562
rect -2 -1598 455 -1568
rect 442 -1603 455 -1598
rect 445 -1608 455 -1603
rect 507 -1608 517 -1556
<< via1 >>
rect 454 508 506 560
rect 197 176 249 228
rect 399 100 451 300
rect 276 10 328 62
rect 116 -154 168 -102
rect -49 -393 3 -193
rect 195 -322 252 -267
rect 441 -323 497 -267
rect -50 -885 2 -685
rect 193 -822 251 -764
rect 440 -818 496 -762
rect 116 -975 168 -923
rect 274 -1139 326 -1087
rect 193 -1305 251 -1247
rect 397 -1377 449 -1177
rect 455 -1608 507 -1556
<< metal2 >>
rect 452 562 508 572
rect 452 496 508 506
rect -42 419 451 461
rect -42 -183 -6 419
rect 399 300 451 419
rect 195 230 251 240
rect 195 164 251 174
rect 399 90 451 100
rect 276 62 328 72
rect 276 -32 328 10
rect 115 -84 328 -32
rect 115 -102 169 -84
rect 115 -154 116 -102
rect 168 -154 169 -102
rect 116 -164 168 -154
rect -49 -193 3 -183
rect 194 -266 252 -256
rect 194 -334 252 -324
rect 441 -267 497 -257
rect 441 -333 497 -323
rect -49 -403 3 -393
rect -42 -675 -6 -403
rect -50 -685 2 -675
rect 193 -764 251 -754
rect 193 -832 251 -822
rect 440 -762 496 -752
rect 440 -828 496 -818
rect -50 -895 2 -885
rect -42 -1481 -6 -895
rect 116 -923 168 -913
rect 116 -1002 168 -975
rect 116 -1048 326 -1002
rect 274 -1087 326 -1048
rect 274 -1149 326 -1139
rect 397 -1177 449 -1167
rect 193 -1247 251 -1237
rect 193 -1315 251 -1305
rect 449 -1377 450 -1316
rect 397 -1481 450 -1377
rect -42 -1516 450 -1481
rect 453 -1554 509 -1544
rect 453 -1620 509 -1610
<< via2 >>
rect 452 560 508 562
rect 452 508 454 560
rect 454 508 506 560
rect 506 508 508 560
rect 452 506 508 508
rect 195 228 251 230
rect 195 176 197 228
rect 197 176 249 228
rect 249 176 251 228
rect 195 174 251 176
rect 194 -267 252 -266
rect 194 -322 195 -267
rect 195 -322 252 -267
rect 194 -324 252 -322
rect 441 -323 497 -267
rect 193 -822 251 -764
rect 440 -818 496 -762
rect 193 -1305 251 -1247
rect 453 -1556 509 -1554
rect 453 -1608 455 -1556
rect 455 -1608 507 -1556
rect 507 -1608 509 -1556
rect 453 -1610 509 -1608
<< metal3 >>
rect 442 562 518 567
rect 442 506 452 562
rect 508 506 518 562
rect 442 501 518 506
rect 185 230 261 235
rect 185 174 195 230
rect 251 174 261 230
rect 185 169 261 174
rect 193 -261 254 169
rect 184 -266 262 -261
rect 453 -262 513 501
rect 184 -324 194 -266
rect 252 -324 262 -266
rect 184 -329 262 -324
rect 431 -267 513 -262
rect 431 -323 441 -267
rect 497 -323 513 -267
rect 431 -328 513 -323
rect 193 -759 254 -329
rect 453 -757 513 -328
rect 183 -764 261 -759
rect 183 -822 193 -764
rect 251 -822 261 -764
rect 183 -827 261 -822
rect 430 -762 513 -757
rect 430 -818 440 -762
rect 496 -818 513 -762
rect 430 -823 513 -818
rect 193 -1242 254 -827
rect 183 -1247 261 -1242
rect 183 -1305 193 -1247
rect 251 -1305 261 -1247
rect 183 -1310 261 -1305
rect 453 -1549 513 -823
rect 443 -1554 519 -1549
rect 443 -1610 453 -1554
rect 509 -1610 519 -1554
rect 443 -1615 519 -1610
use sky130_fd_pr__pfet_01v8_2XU92K  sky130_fd_pr__pfet_01v8_2XU92K_0
timestamp 1729240572
transform 1 0 424 0 1 -785
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU92K  sky130_fd_pr__pfet_01v8_2XU92K_1
timestamp 1729240572
transform 1 0 425 0 1 -293
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU92K  sky130_fd_pr__pfet_01v8_2XU92K_2
timestamp 1729240572
transform 1 0 425 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU92K  sky130_fd_pr__pfet_01v8_2XU92K_3
timestamp 1729240572
transform 1 0 21 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU92K  sky130_fd_pr__pfet_01v8_2XU92K_4
timestamp 1729240572
transform 1 0 21 0 1 -293
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU92K  sky130_fd_pr__pfet_01v8_2XU92K_5
timestamp 1729240572
transform 1 0 20 0 1 -785
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU92K  sky130_fd_pr__pfet_01v8_2XU92K_6
timestamp 1729240572
transform 1 0 19 0 1 -1277
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU92K  sky130_fd_pr__pfet_01v8_2XU92K_7
timestamp 1729240572
transform 1 0 423 0 1 -1277
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_0
timestamp 1729240572
transform 1 0 221 0 1 -1277
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_1
timestamp 1729240572
transform 1 0 223 0 1 200
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_2
timestamp 1729240572
transform 1 0 223 0 1 -293
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_3
timestamp 1729240572
transform 1 0 222 0 1 -785
box -223 -200 223 200
<< labels >>
flabel viali 132 624 132 624 0 FreeSans 320 0 0 0 VDD
port 1 nsew
flabel metal2 112 442 112 442 0 FreeSans 320 0 0 0 D6
port 3 nsew
flabel metal3 221 -107 221 -106 0 FreeSans 320 0 0 0 D5
port 11 nsew
flabel metal3 481 446 481 446 0 FreeSans 320 0 0 0 OUT
port 15 nsew
flabel metal1 300 -993 300 -993 0 FreeSans 320 0 0 0 VIP
port 23 nsew
flabel metal2 298 -11 298 -11 0 FreeSans 320 0 0 0 VIN
port 27 nsew
<< end >>
