magic
tech sky130A
magscale 1 2
timestamp 1729440784
<< viali >>
rect 2410 2819 2462 2871
rect 2409 2685 2461 2737
rect 2160 1759 2240 1853
rect 2299 1775 2333 1842
rect 2428 1425 2480 1477
rect 1743 1139 1781 1175
<< metal1 >>
rect 604 2931 2676 2989
rect 604 2842 662 2931
rect 2410 2886 2462 2931
rect 2397 2871 2475 2886
rect 2397 2819 2410 2871
rect 2462 2819 2475 2871
rect 2397 2808 2475 2819
rect 2396 2737 2474 2752
rect 2144 2655 2154 2707
rect 2206 2655 2216 2707
rect 2396 2685 2409 2737
rect 2461 2685 2474 2737
rect 2396 2674 2474 2685
rect 2407 2644 2463 2674
rect 2407 2609 2540 2644
rect 2227 2524 2237 2576
rect 2289 2524 2299 2576
rect 972 2204 1188 2257
rect 620 2055 1152 2090
rect 620 2054 704 2055
rect 2154 1853 2246 1865
rect 2293 1853 2339 1854
rect 2154 1759 2160 1853
rect 2240 1842 2339 1853
rect 2240 1775 2299 1842
rect 2333 1775 2339 1842
rect 2240 1763 2339 1775
rect 2240 1759 2246 1763
rect 2154 1747 2246 1759
rect 2489 1724 2539 2609
rect 2618 2508 2676 2931
rect 2622 2430 2676 2508
rect 2618 2394 2676 2430
rect 2617 2346 2931 2394
rect 2490 1680 2991 1724
rect 2399 1590 2409 1642
rect 2461 1641 2672 1642
rect 2461 1591 2945 1641
rect 2461 1590 2672 1591
rect 1686 1423 1722 1496
rect 2415 1477 2493 1492
rect 2415 1425 2428 1477
rect 2480 1425 2493 1477
rect 1686 1392 1783 1423
rect 2415 1413 2493 1425
rect 1743 1187 1781 1392
rect 2428 1195 2480 1413
rect 1731 1181 1783 1187
rect 1783 1133 1793 1181
rect 2428 1143 2552 1195
rect 1731 1123 1783 1129
rect 1214 1055 1248 1056
rect 2400 1055 2410 1062
rect 1213 1018 2410 1055
rect 1214 817 1248 1018
rect 2086 818 2120 1018
rect 2400 1010 2410 1018
rect 2462 1010 2472 1062
rect 2271 980 2323 986
rect 2271 465 2323 928
rect 2500 193 2552 1143
rect 2488 135 2498 193
rect 2551 135 2561 193
<< via1 >>
rect 2154 2655 2206 2707
rect 2237 2524 2289 2576
rect 2409 1590 2461 1642
rect 1731 1175 1783 1181
rect 1731 1139 1743 1175
rect 1743 1139 1781 1175
rect 1781 1139 1783 1175
rect 1731 1129 1783 1139
rect 2410 1010 2462 1062
rect 2271 928 2323 980
rect 2498 135 2551 193
<< metal2 >>
rect 2130 2724 2227 2734
rect 2130 2617 2227 2627
rect 2237 2576 2289 2586
rect 2289 2524 2461 2576
rect 2237 2514 2289 2524
rect 972 2261 1028 2271
rect 972 2195 1028 2205
rect 5 1852 61 1862
rect 5 1786 61 1796
rect 2409 1724 2461 2524
rect 2409 1678 2460 1724
rect 2409 1642 2461 1678
rect 2408 1602 2409 1630
rect 2409 1580 2461 1590
rect 1098 1340 1154 1350
rect 610 1285 1098 1340
rect 1154 1285 1155 1340
rect 1098 1274 1154 1284
rect 1725 1129 1731 1181
rect 1783 1129 2323 1181
rect 2271 980 2323 1129
rect 2410 1062 2462 1072
rect 2406 1010 2410 1029
rect 2462 1010 2463 1029
rect 2265 928 2271 980
rect 2323 928 2329 980
rect 2406 611 2463 1010
rect 2539 611 2815 612
rect 2405 610 2815 611
rect 2404 568 2815 610
rect 2119 526 2464 527
rect 1205 473 2464 526
rect 2393 189 2447 473
rect 2497 193 2553 203
rect 2393 137 2497 189
rect 2393 135 2498 137
rect 2551 135 2553 137
rect 2497 127 2553 135
rect 2498 125 2551 127
<< via2 >>
rect 2130 2707 2227 2724
rect 2130 2655 2154 2707
rect 2154 2655 2206 2707
rect 2206 2655 2227 2707
rect 2130 2627 2227 2655
rect 972 2205 1028 2261
rect 5 1796 61 1852
rect 1098 1284 1154 1340
rect 2497 137 2498 193
rect 2498 137 2551 193
rect 2551 137 2553 193
<< metal3 >>
rect 2120 2724 2237 2729
rect 2120 2628 2130 2724
rect 2114 2627 2130 2628
rect 2227 2627 2237 2724
rect 2114 2622 2237 2627
rect 962 2261 1038 2266
rect 962 2205 972 2261
rect 1028 2205 1038 2261
rect 962 2200 1038 2205
rect -5 1852 71 1857
rect -5 1850 5 1852
rect -6 1796 5 1850
rect 61 1796 71 1852
rect -6 1790 71 1796
rect -6 1479 66 1790
rect 971 1479 1031 2200
rect 2114 2184 2224 2622
rect 1720 2124 2224 2184
rect -6 1416 1031 1479
rect 5 1415 1031 1416
rect 971 1414 1031 1415
rect 1088 1342 1164 1345
rect 2771 1342 3072 1343
rect 1088 1340 3072 1342
rect 1088 1284 1098 1340
rect 1154 1284 3072 1340
rect 1088 1280 3072 1284
rect 1088 1279 1164 1280
rect 2771 1279 3072 1280
rect 2487 196 2563 198
rect 2486 193 3339 196
rect 2486 191 2497 193
rect 2484 137 2497 191
rect 2553 137 3339 193
rect 2484 130 3339 137
rect 2484 125 2562 130
rect 2485 122 2562 125
use opamp1  opamp1_1
timestamp 1729429164
transform 1 0 -29 0 1 104
box -178 -106 822 2824
use opamp2  opamp2_0
timestamp 1729431229
transform 1 0 1223 0 1 2207
box -387 -753 1110 642
use opamp3  opamp3_0
timestamp 1729412534
transform 1 0 2821 0 1 1745
box -217 -1748 655 679
use opamp4  opamp4_0
timestamp 1729440198
transform 1 0 1195 0 1 92
box -188 -71 1118 1096
<< labels >>
flabel via1 2262 2547 2262 2547 0 FreeSans 480 0 0 0 VIN
port 6 nsew
flabel viali 2430 2712 2430 2712 0 FreeSans 480 0 0 0 VIP
port 8 nsew
flabel viali 2436 2844 2436 2844 0 FreeSans 320 0 0 0 VDD
port 18 nsew
flabel viali 2451 1451 2451 1451 0 FreeSans 320 0 0 0 OUT
port 22 nsew
flabel via1 2182 2674 2182 2674 0 FreeSans 480 0 0 0 RS
port 10 nsew
flabel viali 2196 1810 2196 1810 0 FreeSans 320 0 0 0 GND
port 24 nsew
<< end >>
