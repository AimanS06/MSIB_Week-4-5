magic
tech sky130A
magscale 1 2
timestamp 1729434446
<< error_s >>
rect 782 2860 930 2894
rect 810 2849 930 2860
rect 964 2849 1000 2875
rect 2328 2849 2359 2875
rect 836 2826 964 2849
rect 836 2823 912 2826
rect 802 2816 912 2823
rect 930 2816 964 2826
rect 1000 2816 1026 2849
rect 802 2815 1026 2816
rect 802 2812 896 2815
rect 802 2796 870 2812
rect 802 2789 828 2796
rect 836 2789 878 2796
rect 836 2762 896 2789
rect 836 2746 870 2762
rect 836 2360 896 2746
rect 2265 2624 2279 2676
rect 2299 2590 2313 2710
rect 2333 2442 2359 2849
rect 2316 2423 2359 2442
rect 2316 2388 2333 2423
rect 828 2326 896 2360
rect 836 2314 870 2326
rect 836 2137 837 2314
rect 870 2137 896 2314
rect 836 2056 896 2137
rect 836 2040 870 2056
rect 214 1851 266 1994
rect 214 1798 267 1851
rect 214 1618 266 1798
rect 836 1652 896 2040
rect 828 1618 896 1652
rect 836 1606 870 1618
rect 836 1457 837 1606
rect 870 1516 896 1606
rect 2131 1585 2168 1635
rect 870 1490 930 1516
rect 964 1490 1000 1516
rect 930 1457 964 1490
rect 1000 1457 1026 1490
rect 836 1456 1026 1457
rect 2334 1456 2359 2423
rect 2370 1456 2387 2388
rect 960 1173 964 1227
rect 988 1173 1000 1199
rect 1014 6 1026 1173
rect 1743 953 1781 989
rect 2334 6 2340 1199
<< nwell >>
rect 0 2928 1003 3100
rect 0 2927 1001 2928
rect 2326 2919 3199 3091
rect 2328 2423 3210 2919
<< viali >>
rect 2227 2824 2279 2876
rect 2227 2624 2279 2676
rect 2259 2401 2311 2453
rect 2259 2295 2311 2347
rect 2131 1585 2168 1635
rect 1743 953 1781 989
<< metal1 >>
rect 816 2931 2676 2989
rect 816 2842 874 2931
rect 2233 2889 2274 2931
rect 2214 2876 2291 2889
rect 2214 2824 2227 2876
rect 2279 2824 2291 2876
rect 2214 2811 2291 2824
rect 2226 2727 2236 2779
rect 2288 2727 2298 2779
rect 2214 2676 2292 2691
rect 2214 2624 2227 2676
rect 2279 2624 2461 2676
rect 2214 2613 2292 2624
rect 2227 2524 2237 2576
rect 2289 2524 2299 2576
rect 2246 2453 2324 2468
rect 2173 2447 2207 2448
rect 2246 2447 2259 2453
rect 2172 2408 2259 2447
rect 972 2204 1188 2257
rect 678 2055 1162 2090
rect 204 1798 214 1851
rect 267 1798 277 1851
rect 2173 1647 2207 2408
rect 2246 2401 2259 2408
rect 2311 2401 2324 2453
rect 2246 2390 2324 2401
rect 2246 2347 2324 2361
rect 2246 2295 2259 2347
rect 2311 2295 2324 2347
rect 2246 2283 2324 2295
rect 2257 2233 2311 2283
rect 2257 2195 2361 2233
rect 2125 1635 2207 1647
rect 2125 1585 2131 1635
rect 2168 1592 2207 1635
rect 2168 1585 2174 1592
rect 2125 1573 2174 1585
rect 1686 1423 1722 1496
rect 1686 1392 1783 1423
rect 1743 1111 1781 1392
rect 1208 1061 1630 1111
rect 1208 816 1254 1061
rect 1620 1059 1630 1061
rect 1682 1061 2125 1111
rect 1682 1059 1692 1061
rect 1743 995 1781 1061
rect 1731 989 1793 995
rect 1731 953 1743 989
rect 1781 953 1793 989
rect 1731 947 1793 953
rect 2081 834 2124 1061
rect 2306 919 2360 2195
rect 2408 1724 2460 2624
rect 2618 2347 2676 2931
rect 2408 1680 2688 1724
rect 2399 1590 2409 1642
rect 2461 1590 2672 1642
rect 1621 167 1631 219
rect 1683 167 1693 219
<< via1 >>
rect 2236 2727 2288 2779
rect 2237 2524 2289 2576
rect 214 1798 267 1851
rect 1630 1059 1682 1111
rect 2409 1590 2461 1642
rect 1631 167 1683 219
<< metal2 >>
rect 2236 2779 2288 2789
rect 2173 2736 2236 2767
rect 972 2261 1028 2271
rect 972 2195 1028 2205
rect 2173 2177 2206 2736
rect 2236 2717 2288 2727
rect 2237 2576 2289 2586
rect 2289 2524 2461 2576
rect 2237 2514 2289 2524
rect 1976 2131 2207 2177
rect 213 1852 269 1862
rect 213 1786 269 1796
rect 2409 1642 2461 2524
rect 2409 1580 2461 1590
rect 1098 1340 1154 1350
rect 817 1285 1098 1340
rect 1154 1285 1155 1340
rect 1098 1274 1154 1284
rect 1628 1113 1684 1123
rect 1628 1047 1684 1057
rect 2305 926 2361 936
rect 2305 860 2361 870
rect 1629 221 1685 231
rect 1629 155 1685 165
<< via2 >>
rect 972 2205 1028 2261
rect 213 1851 269 1852
rect 213 1798 214 1851
rect 214 1798 267 1851
rect 267 1798 269 1851
rect 213 1796 269 1798
rect 1098 1284 1154 1340
rect 1628 1111 1684 1113
rect 1628 1059 1630 1111
rect 1630 1059 1682 1111
rect 1682 1059 1684 1111
rect 1628 1057 1684 1059
rect 2305 870 2361 926
rect 1629 219 1685 221
rect 1629 167 1631 219
rect 1631 167 1683 219
rect 1683 167 1685 219
rect 1629 165 1685 167
<< metal3 >>
rect 962 2261 1038 2266
rect 962 2205 972 2261
rect 1028 2205 1038 2261
rect 962 2200 1038 2205
rect 203 1852 279 1857
rect 203 1796 213 1852
rect 269 1796 279 1852
rect 203 1791 279 1796
rect 214 1479 274 1791
rect 971 1479 1031 2200
rect 214 1415 1031 1479
rect 971 1414 1031 1415
rect 1088 1342 1164 1345
rect 1088 1340 2806 1342
rect 1088 1284 1098 1340
rect 1154 1284 2806 1340
rect 1088 1280 2806 1284
rect 1088 1279 1164 1280
rect 1618 1113 1694 1118
rect 1618 1057 1628 1113
rect 1684 1057 1694 1113
rect 1618 1052 1694 1057
rect 1626 226 1688 1052
rect 2295 926 2371 931
rect 2295 870 2305 926
rect 2361 870 2371 926
rect 2295 865 2371 870
rect 1619 221 1695 226
rect 1619 165 1629 221
rect 1685 165 1695 221
rect 1619 160 1695 165
rect 2295 196 2369 865
rect 1627 82 1687 160
rect 2295 132 3070 196
rect 2295 82 2369 132
rect 1627 46 2369 82
rect 1628 40 2369 46
rect 1628 22 2368 40
use opamp1  opamp1_0
timestamp 1729429164
transform 1 0 178 0 1 106
box -178 -106 822 2824
use opamp2  opamp2_0
timestamp 1729431229
transform 1 0 1223 0 1 2207
box -387 -753 1110 642
use opamp3  opamp3_0
timestamp 1729412534
transform 1 0 2551 0 1 1745
box -217 -1748 655 679
use opamp4  opamp4_0
timestamp 1729434446
transform 1 0 1202 0 1 77
box -188 -71 1118 1096
<< labels >>
flabel viali 2284 2320 2284 2320 0 FreeSans 480 0 0 0 OUT
port 2 nsew
flabel viali 2284 2418 2284 2418 0 FreeSans 480 0 0 0 GND
port 4 nsew
flabel via1 2262 2547 2262 2547 0 FreeSans 480 0 0 0 VIN
port 6 nsew
flabel viali 2248 2651 2248 2651 0 FreeSans 480 0 0 0 VIP
port 8 nsew
flabel via1 2264 2746 2264 2746 0 FreeSans 480 0 0 0 RS
port 10 nsew
flabel viali 2251 2853 2251 2853 0 FreeSans 480 0 0 0 VDD
port 12 nsew
<< end >>
